module register_file(
elk,
nrst,
rd_addrA, rd_addrB, wr_addr, wr_en,
wr_data, rd_dataA, rd_dataB
);
