module module_name ();

endmodule //
